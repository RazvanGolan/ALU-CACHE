library verilog;
use verilog.vl_types.all;
entity ALU_tb is
    generic(
        CLK_PERIOD      : integer := 100
    );
end ALU_tb;
